class miim_agent extends uvm_agent;
	`uvm_component_utils(miim_agent)
	`NEW_COMP
endclass
