typedef uvm_sequencer#(eth_frame) rx_sqr;
