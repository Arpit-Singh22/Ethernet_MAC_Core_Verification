class tx_agent extends uvm_agent;
	`uvm_component_utils(tx_agent)
	`NEW_COMP
endclass
