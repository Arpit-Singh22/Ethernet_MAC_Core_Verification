typedef uvm_sequencer#(wb_tx) proc_sqr;
